`timescale 1ns / 1ps

module tb_sr_latch(

    );
    
reg S,R;
wire Q, Q_bar;


sr_latch uut(S,R,Q,Q_bar);

initial 
    begin
    S=0;  
    R=1;
    #10
    S=1;  
    R=1;
    #10
    S=1;  
    R=0;
    #10
    S=1;  
    R=1;
    #10
    S=0;  
    R=0;
    #10
  $finish;
  end

endmodule