`timescale 1ns / 1ps

module tb_mux_4x1_gates();

reg I0, I1, I2, I3, S0, S1;
wire Y;

mux_4x1_gates uut(I0, I1, I2, I3, S0, S1, Y);

initial begin
    // S1=0, S0=0
    S1=0; S0=0;
    I0=0; I1=0; I2=0; I3=0; #10;
    I0=0; I1=0; I2=0; I3=1; #10;
    I0=0; I1=0; I2=1; I3=0; #10;
    I0=0; I1=0; I2=1; I3=1; #10;
    I0=0; I1=1; I2=0; I3=0; #10;
    I0=0; I1=1; I2=0; I3=1; #10;
    I0=0; I1=1; I2=1; I3=0; #10;
    I0=0; I1=1; I2=1; I3=1; #10;
    I0=1; I1=0; I2=0; I3=0; #10;
    I0=1; I1=0; I2=0; I3=1; #10;
    I0=1; I1=0; I2=1; I3=0; #10;
    I0=1; I1=0; I2=1; I3=1; #10;
    I0=1; I1=1; I2=0; I3=0; #10;
    I0=1; I1=1; I2=0; I3=1; #10;
    I0=1; I1=1; I2=1; I3=0; #10;
    I0=1; I1=1; I2=1; I3=1; #10;

    // S1=0, S0=1
    S1=0; S0=1;
    I0=0; I1=0; I2=0; I3=0; #10;
    I0=0; I1=0; I2=0; I3=1; #10;
    I0=0; I1=0; I2=1; I3=0; #10;
    I0=0; I1=0; I2=1; I3=1; #10;
    I0=0; I1=1; I2=0; I3=0; #10;
    I0=0; I1=1; I2=0; I3=1; #10;
    I0=0; I1=1; I2=1; I3=0; #10;
    I0=0; I1=1; I2=1; I3=1; #10;
    I0=1; I1=0; I2=0; I3=0; #10;
    I0=1; I1=0; I2=0; I3=1; #10;
    I0=1; I1=0; I2=1; I3=0; #10;
    I0=1; I1=0; I2=1; I3=1; #10;
    I0=1; I1=1; I2=0; I3=0; #10;
    I0=1; I1=1; I2=0; I3=1; #10;
    I0=1; I1=1; I2=1; I3=0; #10;
    I0=1; I1=1; I2=1; I3=1; #10;

    // S1=1, S0=0
    S1=1; S0=0;
    I0=0; I1=0; I2=0; I3=0; #10;
    I0=0; I1=0; I2=0; I3=1; #10;
    I0=0; I1=0; I2=1; I3=0; #10;
    I0=0; I1=0; I2=1; I3=1; #10;
    I0=0; I1=1; I2=0; I3=0; #10;
    I0=0; I1=1; I2=0; I3=1; #10;
    I0=0; I1=1; I2=1; I3=0; #10;
    I0=0; I1=1; I2=1; I3=1; #10;
    I0=1; I1=0; I2=0; I3=0; #10;
    I0=1; I1=0; I2=0; I3=1; #10;
    I0=1; I1=0; I2=1; I3=0; #10;
    I0=1; I1=0; I2=1; I3=1; #10;
    I0=1; I1=1; I2=0; I3=0; #10;
    I0=1; I1=1; I2=0; I3=1; #10;
    I0=1; I1=1; I2=1; I3=0; #10;
    I0=1; I1=1; I2=1; I3=1; #10;

    // S1=1, S0=1
    S1=1; S0=1;
    I0=0; I1=0; I2=0; I3=0; #10;
    I0=0; I1=0; I2=0; I3=1; #10;
    I0=0; I1=0; I2=1; I3=0; #10;
    I0=0; I1=0; I2=1; I3=1; #10;
    I0=0; I1=1; I2=0; I3=0; #10;
    I0=0; I1=1; I2=0; I3=1; #10;
    I0=0; I1=1; I2=1; I3=0; #10;
    I0=0; I1=1; I2=1; I3=1; #10;
    I0=1; I1=0; I2=0; I3=0; #10;
    I0=1; I1=0; I2=0; I3=1; #10;
    I0=1; I1=0; I2=1; I3=0; #10;
    I0=1; I1=0; I2=1; I3=1; #10;
    I0=1; I1=1; I2=0; I3=0; #10;
    I0=1; I1=1; I2=0; I3=1; #10;
    I0=1; I1=1; I2=1; I3=0; #10;
    I0=1; I1=1; I2=1; I3=1; #10;

    $finish;
end
endmodule
